module helloworld;
    initial begin
        $display("Hello Verilog");
    end

endmodule